module SDRAM_HY57V641620(
	
);

endmodule
